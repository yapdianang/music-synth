// How to use:					
// 1. Edit the songs on the Enter Song sheet.					
// 2. Select this whole worksheet, copy it, and paste it into a new file.					
// 3. Save the file as song_rom.v.					
					
module song_rom (					
	input clk,				
	input [8:0] addr,				
	output reg [15:0] dout				
);					
					 
	wire [15:0] memory [511:0];				
					
	always @(posedge clk)				 
		dout = memory[addr];			 

assign memory[	  0	] =	{1'b0, 6'd28, 6'd10,  3'b0};	// Note: 3C
assign memory[	  1	] =	{1'b0, 6'd25, 6'd10,  3'b0};	// Note: 3A
assign memory[	  2	] =	{1'b0, 6'd23, 6'd10,  3'b0};	// Note: 2G
assign memory[	  3	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	  4	] =	{1'b0, 6'd28, 6'd10,  3'b0};	// Note: 3C
assign memory[	  5	] =	{1'b0, 6'd25, 6'd10,  3'b0};	// Note: 3A
assign memory[	  6	] =	{1'b0, 6'd23, 6'd10,  3'b0};	// Note: 2G
assign memory[	  7	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	  8	] =	{1'b0, 6'd28, 6'd10,  3'b0};	// Note: 3C
assign memory[	  9	] =	{1'b0, 6'd25, 6'd10,  3'b0};	// Note: 3A
assign memory[	 10	] =	{1'b0, 6'd23, 6'd10,  3'b0};	// Note: 2G
assign memory[	 11	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 12	] =	{1'b0, 6'd28, 6'd22,  3'b0};	// Note: 3C
assign memory[	 13	] =	{1'b0, 6'd25, 6'd22,  3'b0};	// Note: 3A
assign memory[	 14	] =	{1'b0, 6'd23, 6'd22,  3'b0};	// Note: 2G
assign memory[	 15	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 16	] =	{1'b0, 6'd28, 6'd22,  3'b0};	// Note: 3C
assign memory[	 17	] =	{1'b0, 6'd25, 6'd22,  3'b0};	// Note: 3A
assign memory[	 18	] =	{1'b0, 6'd23, 6'd22,  3'b0};	// Note: 2G
assign memory[	 19	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 20	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 21	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 22	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 23	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 24	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 25	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 26	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 27	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 28	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 29	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 30	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 31	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 32	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 33	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 34	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 35	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 36	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 37	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 38	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 39	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 40	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 41	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 42	] =	{1'b0, 6'd25, 6'd24,  3'b0};	// Note: 3A
assign memory[	 43	] =	{1'b0, 6'd22, 6'd24,  3'b0};	// Note: 2F#Gb
assign memory[	 44	] =	{1'b0, 6'd18, 6'd24,  3'b0};	// Note: 2D
assign memory[	 45	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 46	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 47	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 48	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 49	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3G
assign memory[	 50	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 51	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 52	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 53	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3G
assign memory[	 54	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 55	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 56	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 57	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3G
assign memory[	 58	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 59	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 60	] =	{1'b0, 6'd28, 6'd24,  3'b0};	// Note: 3C
assign memory[	 61	] =	{1'b0, 6'd25, 6'd24,  3'b0};	// Note: 3A
assign memory[	 62	] =	{1'b0, 6'd21, 6'd24,  3'b0};	// Note: 2F
assign memory[	 63	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 64	] =	{1'b0, 6'd27, 6'd24,  3'b0};	// Note: 3B
assign memory[	 65	] =	{1'b0, 6'd35, 6'd24,  3'b0};	// Note: 3G
assign memory[	 66	] =	{1'b0, 6'd21, 6'd24,  3'b0};	// Note: 2F
assign memory[	 67	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 68	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 69	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 70	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 71	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 72	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 73	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 74	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 75	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 76	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 77	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 78	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 79	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 80	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 81	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 82	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 83	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 84	] =	{1'b0, 6'd28, 6'd24,  3'b0};	// Note: 3C
assign memory[	 85	] =	{1'b0, 6'd23, 6'd24,  3'b0};	// Note: 2G
assign memory[	 86	] =	{1'b0, 6'd20, 6'd24,  3'b0};	// Note: 2E
assign memory[	 87	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 88	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 89	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 90	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 91	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 92	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 93	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 94	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	 95	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 96	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 97	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	 98	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 99	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	100	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	101	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	102	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	103	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	104	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	105	] =	{1'b0, 6'd20, 6'd48,  3'b0};	// Note: 2E
assign memory[	106	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	107	] =	{1'b1, 6'd0, 6'd48,  3'b0};	// Note: rest
assign memory[	108	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	109	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	110	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	111	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	112	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	113	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	114	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	115	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	116	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	117	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	118	] =	{1'b0, 6'd18, 6'd12,  3'b0};	// Note: 2D
assign memory[	119	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	120	] =	{1'b0, 6'd23, 6'd36,  3'b0};	// Note: 2G
assign memory[	121	] =	{1'b0, 6'd20, 6'd36,  3'b0};	// Note: 2E
assign memory[	122	] =	{1'b1, 6'd0, 6'd36,  3'b0};	// Note: rest
assign memory[	123	] =	{1'b0, 6'd16, 6'd24,  3'b0};	// Note: 2C
assign memory[	124	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	125	] =	{1'b0, 6'd25, 6'd64,  3'b0};	// Note: 3A
assign memory[	126	] =	{1'b0, 6'd21, 6'd64,  3'b0};	// Note: 2F
assign memory[	127	] =	{1'b1, 6'd0, 6'd64,  3'b0};	// Note: rest
assign memory[	128	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	129	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	130	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	131	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	132	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	133	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	134	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	135	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	136	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	137	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	138	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	139	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	140	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	141	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	142	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	143	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	144	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	145	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	146	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	147	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	148	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	149	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	150	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	151	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	152	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	153	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	154	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	155	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	156	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	157	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	158	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	159	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	160	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	161	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	162	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	163	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	164	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	165	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	166	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	167	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	168	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	169	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	170	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	171	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	172	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	173	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	174	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	175	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	176	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	177	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	178	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	179	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	180	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	181	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	182	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	183	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	184	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	185	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	186	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	187	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	188	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	189	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	190	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	191	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	192	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	193	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	194	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	195	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	196	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	197	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	198	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	199	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	200	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	201	] =	{1'b0, 6'd47, 6'd48,  3'b0};	// Note: 4G
assign memory[	202	] =	{1'b1, 6'd0, 6'd48,  3'b0};	// Note: rest
assign memory[	203	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	204	] =	{1'b0, 6'd40, 6'd48,  3'b0};	// Note: 4C
assign memory[	205	] =	{1'b1, 6'd0, 6'd48,  3'b0};	// Note: rest
assign memory[	206	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	207	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	208	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	209	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	210	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	211	] =	{1'b0, 6'd47, 6'd32,  3'b0};	// Note: 4G
assign memory[	212	] =	{1'b1, 6'd0, 6'd32,  3'b0};	// Note: rest
assign memory[	213	] =	{1'b0, 6'd16, 6'd48,  3'b0}; // Note: 2C
assign memory[	214	] =	{1'b0, 6'd40, 6'd32,  3'b0};	// Note: 4C
assign memory[	215	] =	{1'b1, 6'd0, 6'd32,  3'b0};	// Note: rest
assign memory[	216	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	217	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	218	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	219	] =	{1'b1, 6'd11, 6'd8,  3'b0};	// Note: rest
assign memory[	220	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	221	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	222	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	223	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	224	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	225	] =	{1'b0, 6'd38, 6'd8,  3'b0};	// Note: 4A#Bb
assign memory[	226	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	227	] =	{1'b0, 6'd40, 6'd8,  3'b0};	// Note: 4C
assign memory[	228	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	229	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	230	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	231	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	232	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	233	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	234	] =	{1'b0, 6'd38, 6'd8,  3'b0};	// Note: 4A#Bb
assign memory[	235	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	236	] =	{1'b0, 6'd40, 6'd8,  3'b0};	// Note: 4C
assign memory[	237	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	238	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	239	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	240	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	241	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	242	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	243	] =	{1'b0, 6'd38, 6'd8,  3'b0};	// Note: 4A#Bb
assign memory[	244	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	245	] =	{1'b0, 6'd40, 6'd8,  3'b0};	// Note: 4C
assign memory[	246	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	247	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	248	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	249	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	250	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	251	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	252	] =	{1'b0, 6'd38, 6'd16,  3'b0};	// Note: 4A#Bb
assign memory[	253	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	254	] =	{1'b0, 6'd0, 6'd0,  3'b0};	// Note: rest
assign memory[	255	] =	{1'b0, 6'd0, 6'd0,  3'b0};	// Note: rest
assign memory[	256	] =	{1'b0, 6'd1, 6'd12,  3'b0};	// Note: 1A
assign memory[	257	] =	{1'b1, 6'd2, 6'd12,  3'b0};	// Note: rest
assign memory[	258	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 1A#Bb
assign memory[	259	] =	{1'b1, 6'd3, 6'd12,  3'b0};	// Note: rest
assign memory[	260	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 1B
assign memory[	261	] =	{1'b1, 6'd5, 6'd12,  3'b0};	// Note: rest
assign memory[	262	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 1C#Db
assign memory[	263	] =	{1'b1, 6'd7, 6'd12,  3'b0};	// Note: rest
assign memory[	264	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 1D#Eb
assign memory[	265	] =	{1'b1, 6'd8, 6'd12,  3'b0};	// Note: rest
assign memory[	266	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 1E
assign memory[	267	] =	{1'b1, 6'd10, 6'd12,  3'b0};	// Note: rest
assign memory[	268	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 1F#Gb
assign memory[	269	] =	{1'b1, 6'd12, 6'd12,  3'b0};	// Note: rest
assign memory[	270	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 1G#Ab
assign memory[	271	] =	{1'b1, 6'd14, 6'd12,  3'b0};	// Note: rest
assign memory[	272	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2A#Bb
assign memory[	273	] =	{1'b1, 6'd15, 6'd12,  3'b0};	// Note: rest
assign memory[	274	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2B
assign memory[	275	] =	{1'b1, 6'd16, 6'd12,  3'b0};	// Note: rest
assign memory[	276	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2C
assign memory[	277	] =	{1'b1, 6'd17, 6'd12,  3'b0};	// Note: rest
assign memory[	278	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2C#Db
assign memory[	279	] =	{1'b1, 6'd18, 6'd12,  3'b0};	// Note: rest
assign memory[	280	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2D
assign memory[	281	] =	{1'b1, 6'd19, 6'd12,  3'b0};	// Note: rest
assign memory[	282	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2D#Eb
assign memory[	283	] =	{1'b1, 6'd20, 6'd12,  3'b0};	// Note: rest
assign memory[	284	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2E
assign memory[	285	] =	{1'b1, 6'd21, 6'd12,  3'b0};	// Note: rest
assign memory[	286	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2F
assign memory[	287	] =	{1'b1, 6'd22, 6'd12,  3'b0};	// Note: rest
assign memory[	288	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	289	] =	{1'b1, 6'd23, 6'd12,  3'b0};	// Note: rest
assign memory[	290	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2G
assign memory[	291	] =	{1'b1, 6'd24, 6'd12,  3'b0};	// Note: rest
assign memory[	292	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 2G#Ab
assign memory[	293	] =	{1'b1, 6'd25, 6'd12,  3'b0};	// Note: rest
assign memory[	294	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3A
assign memory[	295	] =	{1'b1, 6'd26, 6'd12,  3'b0};	// Note: rest
assign memory[	296	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3A#Bb
assign memory[	297	] =	{1'b1, 6'd27, 6'd12,  3'b0};	// Note: rest
assign memory[	298	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3B
assign memory[	299	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	300	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3C
assign memory[	301	] =	{1'b1, 6'd29, 6'd12,  3'b0};	// Note: rest
assign memory[	302	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3C#Db
assign memory[	303	] =	{1'b1, 6'd30, 6'd12,  3'b0};	// Note: rest
assign memory[	304	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3D
assign memory[	305	] =	{1'b1, 6'd31, 6'd12,  3'b0};	// Note: rest
assign memory[	306	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3D#Eb
assign memory[	307	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	308	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	309	] =	{1'b1, 6'd33, 6'd12,  3'b0};	// Note: rest
assign memory[	310	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3F
assign memory[	311	] =	{1'b1, 6'd34, 6'd12,  3'b0};	// Note: rest
assign memory[	312	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3F#Gb
assign memory[	313	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	314	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	315	] =	{1'b1, 6'd36, 6'd12,  3'b0};	// Note: rest
assign memory[	316	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G#Ab
assign memory[	317	] =	{1'b1, 6'd37, 6'd12,  3'b0};	// Note: rest
assign memory[	318	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4A
assign memory[	319	] =	{1'b1, 6'd38, 6'd12,  3'b0};	// Note: rest
assign memory[	320	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4A#Bb
assign memory[	321	] =	{1'b1, 6'd39, 6'd12,  3'b0};	// Note: rest
assign memory[	322	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4B
assign memory[	323	] =	{1'b1, 6'd40, 6'd12,  3'b0};	// Note: rest
assign memory[	324	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4C
assign memory[	325	] =	{1'b1, 6'd41, 6'd12,  3'b0};	// Note: rest
assign memory[	326	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4C#Db
assign memory[	327	] =	{1'b1, 6'd42, 6'd12,  3'b0};	// Note: rest
assign memory[	328	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4D
assign memory[	329	] =	{1'b1, 6'd43, 6'd12,  3'b0};	// Note: rest
assign memory[	330	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4D#Eb
assign memory[	331	] =	{1'b1, 6'd44, 6'd12,  3'b0};	// Note: rest
assign memory[	332	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4E
assign memory[	333	] =	{1'b1, 6'd45, 6'd12,  3'b0};	// Note: rest
assign memory[	334	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4F
assign memory[	335	] =	{1'b1, 6'd46, 6'd12,  3'b0};	// Note: rest
assign memory[	336	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4F#Gb
assign memory[	337	] =	{1'b1, 6'd47, 6'd12,  3'b0};	// Note: rest
assign memory[	338	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4G
assign memory[	339	] =	{1'b1, 6'd48, 6'd12,  3'b0};	// Note: rest
assign memory[	340	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 4G#Ab
assign memory[	341	] =	{1'b1, 6'd49, 6'd12,  3'b0};	// Note: rest
assign memory[	342	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5A
assign memory[	343	] =	{1'b1, 6'd50, 6'd12,  3'b0};	// Note: rest
assign memory[	344	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5A#Bb
assign memory[	345	] =	{1'b1, 6'd51, 6'd12,  3'b0};	// Note: rest
assign memory[	346	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5B
assign memory[	347	] =	{1'b1, 6'd52, 6'd12,  3'b0};	// Note: rest
assign memory[	348	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5C
assign memory[	349	] =	{1'b1, 6'd53, 6'd12,  3'b0};	// Note: rest
assign memory[	350	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5C#Db
assign memory[	351	] =	{1'b1, 6'd54, 6'd12,  3'b0};	// Note: rest
assign memory[	352	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5D
assign memory[	353	] =	{1'b1, 6'd55, 6'd12,  3'b0};	// Note: rest
assign memory[	354	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5D#Eb
assign memory[	355	] =	{1'b1, 6'd56, 6'd12,  3'b0};	// Note: rest
assign memory[	356	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5E
assign memory[	357	] =	{1'b1, 6'd57, 6'd12,  3'b0};	// Note: rest
assign memory[	358	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5F
assign memory[	359	] =	{1'b1, 6'd58, 6'd12,  3'b0};	// Note: rest
assign memory[	360	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5F#Gb
assign memory[	361	] =	{1'b1, 6'd59, 6'd12,  3'b0};	// Note: rest
assign memory[	362	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5G
assign memory[	363	] =	{1'b1, 6'd60, 6'd12,  3'b0};	// Note: rest
assign memory[	364	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 5G#Ab
assign memory[	365	] =	{1'b1, 6'd61, 6'd12,  3'b0};	// Note: rest
assign memory[	366	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 6A
assign memory[	367	] =	{1'b1, 6'd62, 6'd12,  3'b0};	// Note: rest
assign memory[	368	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 6A#Bb
assign memory[	369	] =	{1'b1, 6'd63, 6'd12,  3'b0};	// Note: rest
assign memory[	370	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 6B
assign memory[	371	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	372	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	373	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	374	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	375	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	376	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	377	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	378	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	379	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	380	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	381	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	382	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	383	] =	{1'b1, 6'd28, 6'd4,  3'b0};	// Note: rest
assign memory[	384	] =	{1'b0, 6'd32, 6'd12,  3'b0};	// Note: 3C
assign memory[	385	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3E
assign memory[	386	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	387	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	388	] =	{1'b0, 6'd32, 6'd12,  3'b0};	// Note: 3C
assign memory[	389	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3E
assign memory[	390	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	391	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	392	] =	{1'b0, 6'd32, 6'd12,  3'b0};	// Note: 3C
assign memory[	393	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3E
assign memory[	394	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	395	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	396	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	397	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	398	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	399	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	400	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	401	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	402	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	403	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	404	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	405	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	406	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	407	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	408	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	409	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	410	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	411	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	412	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	413	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	414	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	415	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	416	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	417	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	418	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	419	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	420	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	421	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	422	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	423	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	424	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	425	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	426	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	427	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	428	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	429	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	430	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	431	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	432	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	433	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	434	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	435	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	436	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	437	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	438	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	439	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	440	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	441	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	442	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	443	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	444	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	445	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	446	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	447	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	448	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	449	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	450	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	451	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	452	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	453	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	454	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	455	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	456	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	457	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	458	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	459	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	460	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	461	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	462	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	463	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	464	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	465	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	466	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	467	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	468	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	469	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	470	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	471	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	472	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	473	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	474	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	475	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	476	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	477	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	478	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	479	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	480	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	481	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	482	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	483	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	484	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	485	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	486	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	487	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	488	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	489	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	490	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	491	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	492	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	493	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	494	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	495	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	496	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	497	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	498	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	499	] =	{1'b1, 6'd28, 6'd12,  3'b0};	// Note: rest
assign memory[	500	] =	{1'b0, 6'd0, 6'd48,  3'b0};	// Note: 3C
assign memory[	501	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	502	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	503	] =	{1'b1, 6'd35, 6'd12,  3'b0};	// Note: rest
assign memory[	504	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3G
assign memory[	505	] =	{1'b1, 6'd32, 6'd12,  3'b0};	// Note: rest
assign memory[	506	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: 3E
assign memory[	507	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	508	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	509	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	510	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
assign memory[	511	] =	{1'b1, 6'd0, 6'd4,  3'b0};	// Note: rest
					
endmodule					
					
					
					
					
					
					
					
					
					
					
					
