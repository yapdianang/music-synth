`define NORMAL 3'b000
`define ADD1 3'b001
`define ADD2 3'b010
`define ADD3 3'b011
`define VIOLIN 3'b100
`define CLARINET 3'b101
`define TRUMPET 3'b110
`define CUSTOM 3'b111


module  note_player #(parameter INSTRUMENT = 3'b000)(
    input clk,
    input reset,
    input play_enable,  // When high we play, when low we don't.
    input [5:0] note_to_load,  // The note to play
    input [5:0] duration_to_load,  // The duration of the note to play
    input load_new_note,  // Tells us when we have a new note to load
    output done_with_note,  // When we are done with the note this stays high.
    input beat,  // This is our 1/48th second beat
    input generate_next_sample,  // Tells us when the codec wants a new sample
    output [15:0] sample_out,  // Our sample output
    output new_sample_ready  // Tells the codec when we've got a sample
);

wire [19:0] fr_out, step_size;

wire release_note;
wire rdy_1, rdy_2, rdy_3, rdy_4, rdy_5, rdy_6, rdy_7;
wire [19:0] out_1, out_2, out_3, out_4, out_5, out_6, out_7;
assign step_size = play_enable ? fr_out:20'b0;

countdown_timer ct(
	.clk(clk),
	.reset(reset),
	.playing(play_enable),
	.load_new(load_new_note),
	.duration(duration_to_load),
	.beat(beat),
	.done(done_with_note)
);

frequency_rom fr(
	.clk(clk),
	.addr(note_to_load),
	.dout(fr_out)
);

sine_reader first_harmonic(
	.clk(clk),
	.reset(reset),
	.step_size(step_size),
	.generate_next(generate_next_sample),
	.sample_ready(rdy_1),
	.sample(out_1)
);

sine_reader second_harmonic(
	.clk(clk),
	.reset(reset),
	.step_size(step_size>>1),
	.generate_next(generate_next_sample),
	.sample_ready(rdy_2),
	.sample(out_2)
);

sine_reader third_harmonic(
	.clk(clk),
	.reset(reset),
	.step_size(step_size>>1 + step_size),
	.generate_next(generate_next_sample),
	.sample_ready(rdy_3),
	.sample(out_3)
);

sine_reader forth_harmonic(
	.clk(clk),
	.reset(reset),
	.step_size(step_size>>2),
	.generate_next(generate_next_sample),
	.sample_ready(rdy_4),
	.sample(out_4)
);

sine_reader fifth_harmonic(
	.clk(clk),
	.reset(reset),
	.step_size(step_size>>2 + step_size),
	.generate_next(generate_next_sample),
	.sample_ready(rdy_5),
	.sample(out_5)
);

sine_reader sixth_harmonic(
	.clk(clk),
	.reset(reset),
	.step_size(step_size>>2 + step_size + step_size),
	.generate_next(generate_next_sample),
	.sample_ready(rdy_6),
	.sample(out_6)
);

sine_reader seventh_harmonic(
	.clk(clk),
	.reset(reset),
	.step_size(step_size>>2 + step_size + step_size + step_size),
	.generate_next(generate_next_sample),
	.sample_ready(rdy_7),
	.sample(out_7)
);

reg [16:0] sample_out_reg;

always @(*) begin
	case (INSTRUMENT)
		`NORMAL: begin
			sample_out_reg =  ($signed(out_1) >>> 1);
		end
		`ADD1: begin
			sample_out_reg = (($signed(out_1) >>> 1) + ($signed(out_2) >>> 2));
		end
		`ADD2: begin
			sample_out_reg =  (($signed(out_1) >>> 1) + ($signed(out_2) >>> 2) + ($signed(out_3) >>> 3));
		end
		`ADD3: begin
			sample_out_reg =  (($signed(out_1) >>> 1) + ($signed(out_2) >>> 2) + ($signed(out_3) >>> 3) + ($signed(out_4) >>> 3));
		end
		`VIOLIN: begin
			sample_out_reg =  (($signed(out_1) >>> 1) + ($signed(out_2) >>> 3) + ($signed(out_3) >>> 5) + ($signed(out_4) >>> 7) + ($signed(out_5) >>> 7) + ($signed(out_6) >>> 8) + ($signed(out_7) >>> 9));
		end
		`CLARINET: begin
			sample_out_reg =  (($signed(out_1) >>> 3) + ($signed(out_2) >>> 6) + ($signed(out_3) >>> 3) + ($signed(out_4) >>> 4) + ($signed(out_5) >>> 3) + ($signed(out_6) >>> 4) + ($signed(out_7) >>> 3));
		end
		`TRUMPET: begin
			sample_out_reg =  (($signed(out_1) >>> 4) + ($signed(out_2) >>> 3) + ($signed(out_3) >>> 3) + ($signed(out_4) >>> 3) + ($signed(out_5) >>> 3) + ($signed(out_6) >>> 3) + ($signed(out_7) >>> 4));
		end
		`CUSTOM: begin
			sample_out_reg =  (($signed(out_1) >>> 3) + ($signed(out_2) >>> 2) + ($signed(out_3) >>> 3) + ($signed(out_4) >>> 5) + ($signed(out_5) >>> 5) + ($signed(out_6) >>> 4) + ($signed(out_7) >>> 4));
		end

	endcase
end

assign sample_out = sample_out_reg;

assign new_sample_ready = (rdy_1 & rdy_2 & rdy_3 & rdy_4 & rdy_5 & rdy_6 & rdy_7);

endmodule
