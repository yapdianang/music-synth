`timescale 1ns / 1ps

module one_pulse_kypd(
    );


endmodule
