// How to use:					
// 1. Edit the songs on the Enter Song sheet.					
// 2. Select this whole worksheet, copy it, and paste it into a new file.					
// 3. Save the file as song_rom.v.					
					
module song_rom (					
	input clk,				
	input [8:0] addr,				
	output reg [15:0] dout				
);					
					
	wire [15:0] memory [255:0];				
					
	always @(posedge clk)				
		dout = memory[addr];			
					
assign memory[	  0	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	  1	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	  2	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	  3	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	  4	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	  5	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	  6	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	  7	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	  8	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	  9	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 10	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 11	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 12	] =	{1'b0, 6'd28, 6'd24,  3'b0};	// Note: 3C
assign memory[	 13	] =	{1'b0, 6'd25, 6'd24,  3'b0};	// Note: 3A
assign memory[	 14	] =	{1'b0, 6'd23, 6'd24,  3'b0};	// Note: 2G
assign memory[	 15	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 16	] =	{1'b0, 6'd28, 6'd24,  3'b0};	// Note: 3C
assign memory[	 17	] =	{1'b0, 6'd25, 6'd24,  3'b0};	// Note: 3A
assign memory[	 18	] =	{1'b0, 6'd23, 6'd24,  3'b0};	// Note: 2G
assign memory[	 19	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 20	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 21	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 22	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 23	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 24	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 25	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 26	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 27	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 28	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 29	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 30	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 31	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 32	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 33	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 34	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 35	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 36	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 37	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 38	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 39	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 40	] =	{1'b0, 6'd22, 6'd12,  3'b0};	// Note: 2F#Gb
assign memory[	 41	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 42	] =	{1'b0, 6'd25, 6'd24,  3'b0};	// Note: 3A
assign memory[	 43	] =	{1'b0, 6'd22, 6'd24,  3'b0};	// Note: 2F#Gb
assign memory[	 44	] =	{1'b0, 6'd18, 6'd24,  3'b0};	// Note: 2D
assign memory[	 45	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 46	] =	{1'b0, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 47	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 48	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 49	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3G
assign memory[	 50	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 51	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 52	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 53	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3G
assign memory[	 54	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 55	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 56	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 57	] =	{1'b0, 6'd35, 6'd12,  3'b0};	// Note: 3G
assign memory[	 58	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 59	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 60	] =	{1'b0, 6'd28, 6'd24,  3'b0};	// Note: 3C
assign memory[	 61	] =	{1'b0, 6'd25, 6'd24,  3'b0};	// Note: 3A
assign memory[	 62	] =	{1'b0, 6'd21, 6'd24,  3'b0};	// Note: 2F
assign memory[	 63	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 64	] =	{1'b0, 6'd27, 6'd24,  3'b0};	// Note: 3B
assign memory[	 65	] =	{1'b0, 6'd35, 6'd24,  3'b0};	// Note: 3G
assign memory[	 66	] =	{1'b0, 6'd21, 6'd24,  3'b0};	// Note: 2F
assign memory[	 67	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 68	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 69	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 70	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 71	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 72	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 73	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 74	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 75	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 76	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 77	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 78	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 79	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 80	] =	{1'b0, 6'd28, 6'd12,  3'b0};	// Note: 3C
assign memory[	 81	] =	{1'b0, 6'd25, 6'd12,  3'b0};	// Note: 3A
assign memory[	 82	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	 83	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 84	] =	{1'b0, 6'd28, 6'd24,  3'b0};	// Note: 3C
assign memory[	 85	] =	{1'b0, 6'd23, 6'd24,  3'b0};	// Note: 2G
assign memory[	 86	] =	{1'b0, 6'd20, 6'd24,  3'b0};	// Note: 2E
assign memory[	 87	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	 88	] =	{1'b0, 6'd27, 6'd12,  3'b0};	// Note: 3B
assign memory[	 89	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 90	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 91	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 92	] =	{1'b0, 6'd23, 6'd12,  3'b0};	// Note: 2G
assign memory[	 93	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 94	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	 95	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 96	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	 97	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	 98	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	 99	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	100	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	101	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	102	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	103	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	104	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	105	] =	{1'b0, 6'd20, 6'd48,  3'b0};	// Note: 2E
assign memory[	106	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	107	] =	{1'b1, 6'd0, 6'd48,  3'b0};	// Note: rest
assign memory[	108	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	109	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	110	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	111	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	112	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	113	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	114	] =	{1'b0, 6'd20, 6'd12,  3'b0};	// Note: 2E
assign memory[	115	] =	{1'b0, 6'd16, 6'd12,  3'b0};	// Note: 2C
assign memory[	116	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	117	] =	{1'b0, 6'd21, 6'd12,  3'b0};	// Note: 2F
assign memory[	118	] =	{1'b0, 6'd18, 6'd12,  3'b0};	// Note: 2D
assign memory[	119	] =	{1'b1, 6'd0, 6'd12,  3'b0};	// Note: rest
assign memory[	120	] =	{1'b0, 6'd23, 6'd36,  3'b0};	// Note: 2G
assign memory[	121	] =	{1'b0, 6'd20, 6'd36,  3'b0};	// Note: 2E
assign memory[	122	] =	{1'b1, 6'd0, 6'd36,  3'b0};	// Note: rest
assign memory[	123	] =	{1'b0, 6'd16, 6'd24,  3'b0};	// Note: 2C
assign memory[	124	] =	{1'b1, 6'd0, 6'd24,  3'b0};	// Note: rest
assign memory[	125	] =	{1'b0, 6'd25, 6'd64,  3'b0};	// Note: 3A
assign memory[	126	] =	{1'b0, 6'd21, 6'd64,  3'b0};	// Note: 2F
assign memory[	127	] =	{1'b1, 6'd0, 6'd64,  3'b0};	// Note: rest
assign memory[	128	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	129	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	130	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	131	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	132	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	133	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	134	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	135	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	136	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	137	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	138	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	139	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	140	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	141	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	142	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	143	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	144	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	145	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	146	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	147	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	148	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	149	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	150	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	151	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	152	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	153	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	154	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	155	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	156	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	157	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	158	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	159	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	160	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	161	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	162	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	163	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	164	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	165	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	166	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	167	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	168	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	169	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	170	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	171	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	172	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	173	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	174	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	175	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	176	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	177	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	178	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	179	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	180	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	181	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	182	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	183	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	184	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	185	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	186	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	187	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	188	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	189	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	190	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	191	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	192	] =	{1'b0, 6'd47, 6'd16,  3'b0};	// Note: 4G
assign memory[	193	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	194	] =	{1'b0, 6'd40, 6'd16,  3'b0};	// Note: 4C
assign memory[	195	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	196	] =	{1'b0, 6'd44, 6'd8,  3'b0};	// Note: 4E
assign memory[	197	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	198	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	199	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	200	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	201	] =	{1'b0, 6'd47, 6'd48,  3'b0};	// Note: 4G
assign memory[	202	] =	{1'b1, 6'd0, 6'd48,  3'b0};	// Note: rest
assign memory[	203	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	204	] =	{1'b0, 6'd40, 6'd48,  3'b0};	// Note: 4C
assign memory[	205	] =	{1'b1, 6'd0, 6'd48,  3'b0};	// Note: rest
assign memory[	206	] =	{1'b0, 6'd16, 6'd48,  3'b0};	// Note: 2C
assign memory[	207	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	208	] =	{1'b0, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	209	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	210	] =	{1'b0, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	211	] =	{1'b0, 6'd47, 6'd32,  3'b0};	// Note: 4G
assign memory[	212	] =	{1'b0, 6'd0, 6'd32,  3'b0};	// Note: rest
assign memory[	213	] =	{1'b0, 6'd16, 6'd48,  3'b0}; // Note: 2C
assign memory[	214	] =	{1'b0, 6'd40, 6'd32,  3'b0};	// Note: 4C
assign memory[	215	] =	{1'b1, 6'd0, 6'd32,  3'b0};	// Note: rest
assign memory[	216	] =	{1'b0, 6'd43, 6'd8,  3'b0};	// Note: 4D#Eb
assign memory[	217	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	218	] =	{1'b0, 6'd45, 6'd8,  3'b0};	// Note: 4F
assign memory[	219	] =	{1'b1, 6'd11, 6'd8,  3'b0};	// Note: rest
assign memory[	220	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	221	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	222	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	223	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	224	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	225	] =	{1'b0, 6'd38, 6'd8,  3'b0};	// Note: 4A#Bb
assign memory[	226	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	227	] =	{1'b0, 6'd40, 6'd8,  3'b0};	// Note: 4C
assign memory[	228	] =	{1'b0, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	229	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	230	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	231	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	232	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	233	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	234	] =	{1'b0, 6'd38, 6'd8,  3'b0};	// Note: 4A#Bb
assign memory[	235	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	236	] =	{1'b0, 6'd40, 6'd8,  3'b0};	// Note: 4C
assign memory[	237	] =	{1'b0, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	238	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	239	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	240	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	241	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	242	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	243	] =	{1'b0, 6'd38, 6'd8,  3'b0};	// Note: 4A#Bb
assign memory[	244	] =	{1'b1, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	245	] =	{1'b0, 6'd40, 6'd8,  3'b0};	// Note: 4C
assign memory[	246	] =	{1'b0, 6'd0, 6'd8,  3'b0};	// Note: rest
assign memory[	247	] =	{1'b0, 6'd11, 6'd48,  3'b0};	// Note: 1G
assign memory[	248	] =	{1'b0, 6'd43, 6'd16,  3'b0};	// Note: 4D#Eb
assign memory[	249	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	250	] =	{1'b0, 6'd35, 6'd16,  3'b0};	// Note: 3G
assign memory[	251	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest
assign memory[	252	] =	{1'b0, 6'd38, 6'd16,  3'b0};	// Note: 4A#Bb
assign memory[	253	] =	{1'b1, 6'd0, 6'd16,  3'b0};	// Note: rest


	assign memory[	254	] =	{1'b0, 6'd0, 6'd0,  3'b0};	// Note: rest
	assign memory[	255	] =	{1'b0, 6'd0, 6'd0,  3'b0};	// Note: rest
					
endmodule					
					
					
					
					
					
					
					
					
					
					
					
					
